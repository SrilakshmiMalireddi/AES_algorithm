----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    12:45:09 07/09/2015 
-- Design Name: 
-- Module Name:    sbox - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity sbox is
port (a : in std_logic_vector(7 downto 0);
		y : out std_logic_vector(7 downto 0));
end sbox;

architecture Behavioral of sbox is

begin
process(a)	
begin
case a is
			when "00000000"=>y<=x"63";
			when "00000001"=>y<=x"7c";
			when "00000010"=>y<=x"77";
			when "00000011"=>y<=x"7b";
			when "00000100"=>y<=x"f2";
			when "00000101"=>y<=x"6b";
			when "00000110"=>y<=x"6f";
			when "00000111"=>y<=x"c5";
			when "00001000"=>y<=x"30";
			when "00001001"=>y<=x"01";
			when "00001010"=>y<=x"67";
			when "00001011"=>y<=x"2b";
			when "00001100"=>y<=x"fe";
			when "00001101"=>y<=x"d7";
			when "00001110"=>y<=x"ab";
			when "00001111"=>y<=x"76";
			when "00010000"=>y<=x"ca";
			when "00010001"=>y<=x"82";
			when "00010010"=>y<=x"c9";
			when "00010011"=>y<=x"7d";
			when "00010100"=>y<=x"fa";
			when "00010101"=>y<=x"59";
			when "00010110"=>y<=x"47";
			when "00010111"=>y<=x"f0";
			when "00011000"=>y<=x"ad";
			when "00011001"=>y<=x"d4";
			when "00011010"=>y<=x"a2";
			when "00011011"=>y<=x"af";
			when "00011100"=>y<=x"9c";
			when "00011101"=>y<=x"a4";
			when "00011110"=>y<=x"72";
			when "00011111"=>y<=x"c0";
			when "00100000"=>y<=x"b7";
			when "00100001"=>y<=x"fd";
			when "00100010"=>y<=x"93";
			when "00100011"=>y<=x"26";
			when "00100100"=>y<=x"36";
			when "00100101"=>y<=x"3f";
			when "00100110"=>y<=x"f7";
			when "00100111"=>y<=x"cc";
			when "00101000"=>y<=x"34";
			when "00101001"=>y<=x"a5";
			when "00101010"=>y<=x"e5";
			when "00101011"=>y<=x"f1";
			when "00101100"=>y<=x"71";
			when "00101101"=>y<=x"d8";
			when "00101110"=>y<=x"31";
			when "00101111"=>y<=x"15";
			when "00110000"=>y<=x"04";
			when "00110001"=>y<=x"c7";
			when "00110010"=>y<=x"23";
			when "00110011"=>y<=x"c3";
			when "00110100"=>y<=x"18";
			when "00110101"=>y<=x"96";				
			when "00110110"=>y<=x"05";
			when "00110111"=>y<=x"9a";
			when "00111000"=>y<=x"07";
			when "00111001"=>y<=x"12";
			when "00111010"=>y<=x"80";
			when "00111011"=>y<=x"e2";
			when "00111100"=>y<=x"eb";
			when "00111101"=>y<=x"27";
			when "00111110"=>y<=x"b2";
			when "00111111"=>y<=x"75";
			when "01000000"=>y<=x"09";
			when "01000001"=>y<=x"83";
			when "01000010"=>y<=x"2c";
			when "01000011"=>y<=x"1a";
			when "01000100"=>y<=x"1b";
			when "01000101"=>y<=x"6e";
			when "01000110"=>y<=x"5a";
         when "01000111"=>y<=x"a0";
			when "01001000"=>y<=x"52";
			when "01001001"=>y<=x"3b";
			when "01001010"=>y<=x"d6";
			when "01001011"=>y<=x"b3";
			when "01001100"=>y<=x"29";
			when "01001101"=>y<=x"e3";
			when "01001110"=>y<=x"2f";
		   when "01001111"=>y<=x"84";
			when "01010000"=>y<=x"53";
			when "01010001"=>y<=x"d1";
			when "01010010"=>y<=x"00";
			when "01010011"=>y<=x"ed";
			when "01010100"=>y<=x"20";
			when "01010101"=>y<=x"fc";
			when "01010110"=>y<=x"b1";
			when "01010111"=>y<=x"5b";
			when "01011000"=>y<=x"6a";
			when "01011001"=>y<=x"cb";
			when "01011010"=>y<=x"be";
			when "01011011"=>y<=x"39";
			when "01011100"=>y<=x"4a";
			when "01011101"=>y<=x"4c";
			when "01011110"=>y<=x"58";
			when "01011111"=>y<=x"cf";
			when "01100000"=>y<=x"d0";
			when "01100001"=>y<=x"ef";
			when "01100010"=>y<=x"aa";
			when "01100011"=>y<=x"fb";
			when "01100100"=>y<=x"43";
			when "01100101"=>y<=x"4d";
			when "01100110"=>y<=x"33";
			when "01100111"=>y<=x"85";
			when "01101000"=>y<=x"45";
			when "01101001"=>y<=x"f9";
		   when "01101010"=>y<=x"02";
			when "01101011"=>y<=x"7f";
			when "01101100"=>y<=x"50";
			when "01101101"=>y<=x"3c";
			when "01101110"=>y<=x"9f";
			when "01101111"=>y<=x"a8";
			when "01110000"=>y<=x"51";
			when "01110001"=>y<=x"a3";
			when "01110010"=>y<=x"40";
			when "01110011"=>y<=x"8f";
			when "01110100"=>y<=x"92";
			when "01110101"=>y<=x"9d";
			when "01110110"=>y<=x"38";
		   when "01110111"=>y<=x"f5";
			when "01111000"=>y<=x"bc";
			when "01111001"=>y<=x"b6";
			when "01111010"=>y<=x"da";
			when "01111011"=>y<=x"21";
			when "01111100"=>y<=x"10";
			when "01111101"=>y<=x"ff";
			when "01111110"=>y<=x"f3";
			when "01111111"=>y<=x"d2";
			when "10000000"=>y<=x"cd";
			when "10000001"=>y<=x"0c";
			when "10000010"=>y<=x"13";
			when "10000011"=>y<=x"ec";
			when "10000100"=>y<=x"5f";
			when "10000101"=>y<=x"97";
			when "10000110"=>y<=x"44";
			when "10000111"=>y<=x"17";
			when "10001000"=>y<=x"c4";
			when "10001001"=>y<=x"a7";
			when "10001010"=>y<=x"7e";
			when "10001011"=>y<=x"3d";
			when "10001100"=>y<=x"64";
			when "10001101"=>y<=x"5d";
			when "10001110"=>y<=x"19";
			when "10001111"=>y<=x"73";
			when "10010000"=>y<=x"60";
			when "10010001"=>y<=x"81";
			when "10010010"=>y<=x"4f";
			when "10010011"=>y<=x"dc";
			when "10010100"=>y<=x"22";
			when "10010101"=>y<=x"2a";
			when "10010110"=>y<=x"90";
			when "10010111"=>y<=x"88";
			when "10011000"=>y<=x"46";
			when "10011001"=>y<=x"ee";
			when "10011010"=>y<=x"b8";
			when "10011011"=>y<=x"14";
			when "10011100"=>y<=x"de";
			when "10011101"=>y<=x"5e";
			when "10011110"=>y<=x"0b";
			when "10011111"=>y<=x"db";
			when "10100000"=>y<=x"e0";
			when "10100001"=>y<=x"32";
			when "10100010"=>y<=x"3a";
			when "10100011"=>y<=x"0a";
			when "10100100"=>y<=x"49";
			when "10100101"=>y<=x"06";
			when "10100110"=>y<=x"24";
			when "10100111"=>y<=x"5c";
			when "10101000"=>y<=x"c2";
			when "10101001"=>y<=x"d3";
			when "10101010"=>y<=x"ac";
			when "10101011"=>y<=x"62";
			when "10101100"=>y<=x"91";
			when "10101101"=>y<=x"95";
			when "10101110"=>y<=x"e4";
			when "10101111"=>y<=x"79";
			when "10110000"=>y<=x"e7";
			when "10110001"=>y<=x"c8";
			when "10110010"=>y<=x"37";
			when "10110011"=>y<=x"6d";
			when "10110100"=>y<=x"8d";
			when "10110101"=>y<=x"d5";
			when "10110110"=>y<=x"4e";
			when "10110111"=>y<=x"a9";
			when "10111000"=>y<=x"6c";
			when "10111001"=>y<=x"56";
			when "10111010"=>y<=x"f4";
			when "10111011"=>y<=x"ea";
			when "10111100"=>y<=x"65";
			when "10111101"=>y<=x"7a";
			when "10111110"=>y<=x"ae";
			when "10111111"=>y<=x"08";
			when "11000000"=>y<=x"ba";
			when "11000001"=>y<=x"78";
			when "11000010"=>y<=x"25";
			when "11000011"=>y<=x"2e";
			when "11000100"=>y<=x"1c";
			when "11000101"=>y<=x"a6";
			when "11000110"=>y<=x"b4";
			when "11000111"=>y<=x"c6";
			when "11001000"=>y<=x"e8";
			when "11001001"=>y<=x"dd";
			when "11001010"=>y<=x"74";
			when "11001011"=>y<=x"1f";
			when "11001100"=>y<=x"4b";
			when "11001101"=>y<=x"bd";
			when "11001110"=>y<=x"8b";
			when "11001111"=>y<=x"8a";
			when "11010000"=>y<=x"70";
			when "11010001"=>y<=x"3e";
			when "11010010"=>y<=x"b5";
			when "11010011"=>y<=x"66";
			when "11010100"=>y<=x"48";
			when "11010101"=>y<=x"03";
			when "11010110"=>y<=x"f6";
		   when "11010111"=>y<=x"0e";
			when "11011000"=>y<=x"61";
			when "11011001"=>y<=x"35";
			when "11011010"=>y<=x"57";
			when "11011011"=>y<=x"b9";
			when "11011100"=>y<=x"86";
			when "11011101"=>y<=x"c1";
			when "11011110"=>y<=x"1d";
			when "11011111"=>y<=x"9e";
			when "11100000"=>y<=x"e1";
			when "11100001"=>y<=x"f8";
			when "11100010"=>y<=x"98";
			when "11100011"=>y<=x"11";
			when "11100100"=>y<=x"69";
			when "11100101"=>y<=x"d9";
			when "11100110"=>y<=x"8e";
			when "11100111"=>y<=x"94";
			when "11101000"=>y<=x"9b";
			when "11101001"=>y<=x"1e";
			when "11101010"=>y<=x"87";
			when "11101011"=>y<=x"e9";
			when "11101100"=>y<=x"ce";
			when "11101101"=>y<=x"55";
			when "11101110"=>y<=x"28";
			when "11101111"=>y<=x"df";
			when "11110000"=>y<=x"8c";
			when "11110001"=>y<=x"a1";
			when "11110010"=>y<=x"89";
			when "11110011"=>y<=x"0d";
			when "11110100"=>y<=x"bf";
			when "11110101"=>y<=x"e6";
			when "11110110"=>y<=x"42";
			when "11110111"=>y<=x"68";
			when "11111000"=>y<=x"41";
			when "11111001"=>y<=x"99";
			when "11111010"=>y<=x"2d";
			when "11111011"=>y<=x"0f";
			when "11111100"=>y<=x"b0";
			when "11111101"=>y<=x"54";
			when "11111110"=>y<=x"bb";
			when "11111111"=>y<=x"16";
			
			when others=> y <= x"00";


end case;
end process;
end Behavioral;